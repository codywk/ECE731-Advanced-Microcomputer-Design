module QuadratureEncoderTop (
	input clk,
	input reset,
	input A,
	input B,
	
	);
	
	reg[N-1:0] fwd, mp, bck; // these registers will save the values for specific points to keep track of total distance
	
endmodule
