library verilog;
use verilog.vl_types.all;
entity QuadratureEncoderTop_vlg_vec_tst is
end QuadratureEncoderTop_vlg_vec_tst;
