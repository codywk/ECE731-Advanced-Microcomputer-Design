library verilog;
use verilog.vl_types.all;
entity EncoderPulseCounterTop_vlg_vec_tst is
end EncoderPulseCounterTop_vlg_vec_tst;
